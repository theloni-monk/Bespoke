//WRITEME: ReLU