//WRITEME: dual fifo point-wise ultiplication