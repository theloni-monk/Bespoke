//WRITEME: integrationi netowrk