//TODO: Dual-port BRAM based FIFO with byte masking