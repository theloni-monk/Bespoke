//WRITEME: adder tree
`timescale 1ns / 1ps
`default_nettype none // prevents system from inferring an undeclared logic (good practice)

`default_nettype wire