//WRITME: Dual FIFO point-wise addition