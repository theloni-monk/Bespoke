//WRITEME: Dual FIFO point-wise addition