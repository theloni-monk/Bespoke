//TODO: Dual-port BRAM based FIFO that reads only a few at a time but has